`include "parameters.svh"

module sigmoid
  ( input clk
  , input xrst
  , input enable
  , input out_en
  , input signed [DWIDTH-1:0] pixel_in
  , output signed [DWIDTH-1:0] pixel_out
  );

endmodule
