`include "parameters.svh"

module ctrl_core
  ( input   clk
  , input   xrst
  , input   req
  , output  ack
  );

endmodule
