`ifndef __PARAMETERS_SVH_
`define __PARAMETERS_SVH_

`default_nettype wire
`timescale 1 ns / 1 ps

parameter STEP    = 10;
parameter DWIDTH  = 16;
parameter LWIDTH  = 16;

parameter WAVSIZE = 16;

parameter CORE    = 4;
parameter CORELOG = 2;
parameter NETSIZE = 10;

`endif
