`include "parameters.svh"

module extract
  ( input   clk
  , input   xrst
  );

endmodule
